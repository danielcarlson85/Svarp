﻿--Detta är en kommentar

{variabel}"Detta är värdet i variabeln"
(Skriv){variabel}

{nummer}(RäknaUt)"34*44"
(Skriv){nummer}


(Läs)"Vad heter du? "{var1}
(Skriv)="Hej "{var1}
