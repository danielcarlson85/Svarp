﻿--Detta är en kommentar

{variabel5}(Läs)
{variabel6}(Läs)"Vad heter du? "

(SkrivVariabel){variabel6}





{nummers}"1+1"


(SkrivVariabel){nummers}


(Skriv)"hej"
(RäknaUt)"4+4"





(RäknaUtVariable){nummers}

(SkrivVariabel){nummers}




{variabel1}(Läs)"hej"





(SkrivVariabel){nummers}

(RäknaUt)"22+22"

{variabel2}"Detta är värdet i variabeln"
(Skriv){variabel2}

(RäknaUt)"34*44"


(Läs)"Vad heter du? "{var1}
(Skriv)"Hej "{var1}
