﻿(Läs){input1}
{input2}(Läs)

(Skriv){input2}
(Skriv){input1}


{var1}="första variablen från variable"
(Skriv){var1}



(Skriv)="första raden direkt text"
{var6}="yoyo från variable"
(Skriv)={var6}