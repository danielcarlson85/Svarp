﻿{var1}="första variabel"


(Skriv)"hej"

{input1}(Läs)
{input2}(Läs)

(Skriv){input2}


(Skriv){var1}



(Skriv)="första raden direkt text"
{var6}="yoyo från variable"
(Skriv)={var6}