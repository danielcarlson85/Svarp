﻿//Detta är en kommentar

(Läs)"Vad heter du? "{var1}

(Skriv)="Hej "{var1}