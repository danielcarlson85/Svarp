﻿{variable1}(Läs)"Vad heter du?"
(Skriv)"Vad roligt att du är här:"{test}
{variable2}"När är du född?"(Läs)













SWarp is a swedish sharp programming language that is build for fun

To use:

declare variables: use {}
eg

{variableName1}

Usable methods:
	(Skriv)
	(Läs)
