﻿--Detta är en kommentar
{nummers}"45*23"
(RäknaUt){nummers}
(Skriv){nummers}

(RäknaUt)"22+22"

{variabel}"Detta är värdet i variabeln"
(Skriv){variabel}

{nummer}(RäknaUt)"34*44"
(Skriv){nummer}


(Läs)"Vad heter du? "{var1}
(Skriv)="Hej "{var1}
