﻿(Skriv)"första raden"
{var1}"första variablen"
(Skriv){var1}

{variable1}(Läs)
(Skriv)"Vad roligt att du är här:" {variable1}
{variable2}"När är du född?"(Läs)