﻿(Skriv)			"Jag heter johan vad heter du? "
(Läs)           {variabel1}
(Skriv)			"Vad roligt att du är här " {variabel1}