﻿(Läs){input2}"Hej vad heter du? "
{var1}="första variabel"


(Skriv)"hej"

{input1}(Läs)

(Skriv){input1}

(Skriv){input2}
(Skriv){var1}


(Skriv)="första raden direkt text"
{var6}="yoyo från variable"
(Skriv)={var6}