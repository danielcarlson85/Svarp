﻿//Daniel
(Läs)"Vad heter du? "{var1}


//Johan
(Skriv)="Hej "{var1}