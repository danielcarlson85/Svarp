﻿(Skriv)="första raden"
{var1}="första variablen"
(Skriv){var1}

{var6}="yoyo"

(Skriv){var6}