﻿--Detta är en kommentar

{namn}(LäsInklTitel)"Vad heter du? "
{ålder}(LäsInklTitel)"Hur gammal är du?"
(SkrivUtVariabelOchText){namn}"Välkommen "
(SkrivUtVariabelOchText){ålder}"Du är "




{nummers}"variabel tjoho"


(SkrivVariabel){nummers}


(Skriv)"hej"
(RäknaUt)"4+4"





(RäknaUtVariable){nummers}

(SkrivVariabel){nummers}




{variabel1}(Läs)"hej"





{variabel6}"Daniel"
(SkrivVariabelOchText){variabel6}"hej "

(SkrivVariabel){nummers}

(RäknaUt)"22+22"

{variabel2}"Detta är värdet i variabeln"
(Skriv){variabel2}

(RäknaUt)"34*44"


(Läs)"Vad heter du? "{var1}
(Skriv)"Hej "{var1}


--{nummers}(LäsInklTitel)"Räkna ut: "
--(RäknaUtVariabel){nummers}
--(SkrivUtVariabelOchText){nummers}"Detta skrivs ut också"
--(SkrivUtVariabel){nummers}